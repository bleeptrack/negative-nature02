// Blackbox definition for my_logo module
// This file provides the module definition needed for gate-level testing
(* blackbox *) (* keep *)
module my_logo ();
endmodule
